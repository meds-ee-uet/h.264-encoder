module me #
(
    parameter MACRO_DIM,
    parameter SEARCH_DIM
) 
(
    input  logic        rst_n,
    input  logic        clk,
    input  logic        start,
    input  logic [7:0]  pixel_spr_in [0:MACRO_DIM],
    input  logic [7:0]  pixel_cpr_in [0:MACRO_DIM-1],
    output logic        readyi,
    output logic        en_ram,
    output logic        en_cpr,
    output logic        en_spr,
    input  logic        readyo,
    output logic        valido,
    output logic [5:0]  addr,
    output logic [5:0]  amt,
    output logic [5:0]  mv_x,
    output logic [5:0]  mv_y,
    output logic [15:0] min_sad
);

    logic [1:0] sel;

    datapath_me # 
    (
        .MACRO_DIM  ( MACRO_DIM  ),
        .SEARCH_DIM ( SEARCH_DIM )
    )
    ins_datapath_me
    (
        .rst_n              ( rst_n              ),
        .clk                ( clk                ),
        .amt                ( amt                ),
        .addr               ( addr               ),
        .en_spr             ( en_spr             ),
        .en_cpr             ( en_cpr             ),
        .comp_en            ( comp_en            ),
        .sel                ( sel                ),
        .pixel_spr_in       ( pixel_spr_in       ),
        .pixel_cpr_in       ( pixel_cpr_in       ),
        .min_sad            ( min_sad            ),
        .mv_x               ( mv_x               ),
        .mv_y               ( mv_y               )
    );

    controller_me # 
    (
        .MACRO_DIM  ( MACRO_DIM  ),
        .SEARCH_DIM ( SEARCH_DIM )
    )
    ins_controller_me
    (
        .rst_n      ( rst_n     ), 
        .clk        ( clk       ), 
        .start      ( start     ),
        .readyi     ( readyi    ),
        .comp_en    ( comp_en   ),
        .en_cpr     ( en_cpr    ), 
        .en_spr     ( en_spr    ),
        .en_ram     ( en_ram    ),
        .readyo     ( readyo    ),
        .valido     ( valido    ),
        .addr       ( addr      ),
        .amt        ( amt       ),
        .sel        ( sel       )
    );

endmodule